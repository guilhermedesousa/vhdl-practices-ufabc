library verilog;
use verilog.vl_types.all;
entity xor_schematic_vlg_vec_tst is
end xor_schematic_vlg_vec_tst;
