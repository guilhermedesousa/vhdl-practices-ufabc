library verilog;
use verilog.vl_types.all;
entity paridade_herarquico_vlg_vec_tst is
end paridade_herarquico_vlg_vec_tst;
